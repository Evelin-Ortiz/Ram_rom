library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAM is 
port ( 
		 clock    : in  std_logic;
       address  : in  std_logic_vector(7 downto 0);
		 data_in  : in  std_logic_vector(7 downto 0);
		 WE       : in  std_logic;
		 data_out : out std_logic_vector(7 downto 0));
end entity;
 
 architecture RAM128x8 of RAM is
 
 type rw_type is array (128 to 223) of std_logic_vector(7 downto 0);
signal EN : std_logic;
signal RW : rw_type;
 
 BEGin
 enable : process (address)
 begin
 if ((to_integer(unsigned(address)) >= 128) and
     (to_integer(unsigned(address)) <= 223)) then
	  EN <= '1';
	  else
	  EN <= '0';
	  end if;
end process;
	  
 memory : process (clock)
 begin
   if (clock'event and clock='1') then
   if (EN='1' and WE='1') then
   RW(to_integer(unsigned(address))) <= data_in;
   elsif (EN='1' and WE='0') then
   data_out <= RW(to_integer(unsigned(address)));
   end if;
  end if;
end process;
end architecture;
